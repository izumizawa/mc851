module soc (
    input clk, reset
);

endmodule
